parameter SERIAL = 50;
parameter BATCH = 1;
