parameter SERIAL = 47;
parameter BATCH = 1;
