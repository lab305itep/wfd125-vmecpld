parameter SERIAL = 56;
parameter BATCH = 1;
