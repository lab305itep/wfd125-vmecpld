
parameter SERIAL = 1;
parameter BATCH = 1;
